// module intermediate_register(input  logic clk, reset
//                              input  logic input InputRegister,
//                              output logic input OutputRegtister);

//     always_ff @(posedge clk) begin
//         if (reset)
//             OutputRegtister <= 0;
//         else
//             OutputRegtister <= InputRegister;
//     end

// endmodule